----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/21/2020 11:31:12 PM
-- Design Name: 
-- Module Name: cortex_m0_core - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

library xil_defaultlib;
use xil_defaultlib.helper_funcs.all;


entity cortex_m0_core is
    generic (S_PROGRAM_MEMORY_ENDIAN: boolean := FALSE);           -- little endian = 0, big endian = 1
    Port ( 
            HCLK : in std_logic;                        -- Clock
         HRESETn : in std_logic;                        -- Asynchronous reset

            -- AMBA 3 AHB-LITE INTERFACE INPUTS
          HRDATA : in std_logic_vector (31 downto 0);   -- AHB read-data
          HREADY : in std_logic;                        -- AHB stall signal
           HRESP : in std_logic;                        -- AHB error response

            -- INTERRUPT INPUTS
             NMI : in std_logic;
             IRQ : in std_logic_vector (15 downto 0);
            
            -- EVENT INPUT
            RXEV : in std_logic;
            
--            -- Accelerator related signals:
--            invoke_accelerator : in std_logic;

            -- AMBA 3 AHB-LITE INTERFACE OUTPUTS
           HADDR : out std_logic_vector (31 downto 0);  -- AHB transaction address  format [Lower byte-Upper byte | Lower byte-Upper byte]
          HBURST : out std_logic_vector (2 downto 0);   -- AHB burst: tied to single
       HMASTLOCK : out std_logic;                       -- AHB locked transfer (always zero)
           HPROT : out std_logic_vector (3 downto 0);   -- AHB protection: priv; data or inst
           HSIZE : out std_logic_vector (2 downto 0);   -- AHB size: byte, half-word or word
          HTRANS : out std_logic_vector (1 downto 0);   -- AHB transfer: non-sequential only
          HWDATA : out std_logic_vector (31 downto 0);  -- AHB write-data
          HWRITE : out std_logic;                       -- AHB write control
            
            -- STATUS OUPUTS
        LOCKUP   : out std_logic;    
      SLEEPING   : out std_logic;    
   SYSTESETREQ   : out std_logic;    
            
            -- EVENT OUTPUT
          TXEV   : out std_logic
        );
end cortex_m0_core;

architecture Behavioral of cortex_m0_core is

    -- Components
    component registers is
    Port (
        clk : in std_logic;
        reset : in std_logic;
        WE : in std_logic;
        gp_WR_addr: in std_logic_vector(3 downto 0);
        gp_data_in : in std_logic_vector(31 downto 0);
        gp_addrA: in std_logic_vector(3 downto 0);
        gp_addrB: in std_logic_vector(3 downto 0);
        gp_addrC: in std_logic_vector(3 downto 0);
        gp_ram_dataA : out std_logic_vector(31 downto 0);
        gp_ram_dataB : out std_logic_vector(31 downto 0);
        gp_ram_dataC : out std_logic_vector(31 downto 0)
    );
    end component;
    
    component decoder is
    Port ( 
        clk : in std_logic;
        reset : in std_logic;
        instruction : in std_logic_vector (15 downto 0);
        inst32_detected_in_prev_inst : in boolean;
        inst32_detected : out boolean;
        destination_is_PC : out boolean;
        gp_WR_addr : out STD_LOGIC_VECTOR (3 downto 0);
        gp_addrA: out STD_LOGIC_VECTOR (3 downto 0);
        gp_addrB: out STD_LOGIC_VECTOR (3 downto 0);
        gp_addrC : out std_logic_vector (3 downto 0);
        imm8: out STD_LOGIC_VECTOR (7 downto 0);
        LR_PC : out std_logic;
        execution_cmd: out executor_cmds_t;
        access_mem: out boolean;
        use_base_register : out boolean;
        mem_load_size : out mem_op_size_t;
        mem_load_sign_ext : out boolean;
        LDM_STM_access_mem : out boolean;
        access_mem_mode : out access_mem_mode_t;
        cond : out std_logic_vector (3 downto 0);
        prev_inst : out std_logic_vector (15 downto 0)
    );
    end component;
    
    component executor is
        Port (
             clk : in std_logic;
             reset : in std_logic;
             operand_A : in std_logic_vector(31 downto 0);	
             operand_B : in std_logic_vector(31 downto 0);	
             command: in executor_cmds_t;	
             imm8_z_ext : in  std_logic_vector(31 downto 0);
             destination_is_PC : in boolean;
             current_flags : in flag_t;
             access_mem : in boolean;
             gp_data_in_ctrl : in gp_data_in_ctrl_t;
             disable_executor : in boolean;
             SP_main : in std_logic_vector(31 downto 0);
             cmd_out: out executor_cmds_t;
             set_flags : out boolean;
             result : out std_logic_vector(31 downto 0);
             alu_temp_32 : out std_logic;
             overflow_status : out std_logic_vector(2 downto 0);
             WE: out std_logic;
             SP_updated : out boolean
         );
    end component;
    
    component core_state is
        Port (
            clk : in std_logic;
            reset : in std_logic;
--            instruction_size : in boolean;      -- false = 16-bit (2 bytes), true = 32-bit (4 bytes) 
            access_mem : in boolean;
            PC_updated : in boolean;
            cond : in std_logic_vector (3 downto 0);
            current_flags : in flag_t;
            imm8 : in std_logic_vector (7 downto 0);
            imm8_value : in std_logic_vector (7 downto 0);
            imm11_10_downto_8 : in std_logic_vector (2 downto 0);
            imm11_value_10_downto_8 : in std_logic_vector (2 downto 0);
            LR_PC : in std_logic;
            number_of_ones_initial : in  STD_LOGIC_VECTOR (3 downto 0);
            execution_cmd_value : in executor_cmds_t;
            LDM_STM_access_mem : in boolean;
            new_PC : in std_logic_vector (31 downto 0);
            SP_updated : in boolean;
            access_mem_mode : in access_mem_mode_t;
            SP_main_init : in std_logic_vector (31 downto 0);
            PC_init : in std_logic_vector (31 downto 0);
            pos_A_is_multi_cycle : in boolean;
            ldm_hrdata_value : in std_logic_vector (31 downto 0);
--            hrdata_program : in std_logic_vector(31 downto 0);
            inst32_detected_value : in boolean;
            current_instruction_32bit_HI : in std_logic_vector (15 downto 0);
            current_instruction : in std_logic_vector (15 downto 0);
            msr_update_MSP : in boolean;
            msr_update_PSP : in boolean;
            msr_update_PRIMASK : in boolean;   
            msr_update_CONTROL : in boolean;
            new_PRIMASK : std_logic_vector (0 downto 0);
            new_CONTROL : std_logic_vector (1 downto 0);
            new_SP : in std_logic_vector (31 downto 0);
            PC : out std_logic_vector(31 downto 0);
            SP_main : out std_logic_vector (31 downto 0);
            SP_process : out std_logic_vector (31 downto 0);
            PC_decode : out std_logic_vector (31 downto 0);
            PC_execute :  out std_logic_vector (31 downto 0);
            PC_after_execute :  out std_logic_vector (31 downto 0);
            LDM_STM_mem_address_index :  out unsigned (4 downto 0);          
            gp_data_in_ctrl : out gp_data_in_ctrl_t;
            hrdata_ctrl : out hrdata_ctrl_t;
            disable_fetch : out boolean;
            haddr_ctrl : out haddr_ctrl_t; 
            disable_executor : out boolean;
            gp_addrA_executor_ctrl : out boolean;
            LDM_W_STM_R_reg : out std_logic_vector (3 downto 0);
            LDM_STM_capture_base : out boolean;
            HWRITE : out std_logic;
            VT_ctrl : out VT_ctrl_t;
            branch_target_address : out std_logic_vector (31 downto 0);
            branch_target_address_val : out std_logic_vector (31 downto 0);
            SDC_push_read_address : out SDC_push_read_address_t;
            inst32_detected : out boolean;
            Rn : out std_logic_vector (31 downto 28);
            PRIMASK : out std_logic_vector (0 downto 0);
            CONTROL : out std_logic_vector (1 downto 0)
        );
    end component;
    
     component status_flags is
        Port (
            clk : in std_logic;
            reset : in std_logic;
            result : in std_logic_vector(31 downto 0);
            C_in : in std_logic;
            overflow_status : in std_logic_vector(2 downto 0);
            cmd: in executor_cmds_t;
            set_flags : in boolean; 
            msr_flags : in boolean;
            Rn_content : in std_logic_vector(31 downto 28);                 
            flags_o : out flag_t;
            xPSR : out std_logic_vector(31 downto 0)
            );
    end component;
    
    component count_ones is
        Port ( byte_in : in STD_LOGIC_VECTOR (7 downto 0);
               ones : out STD_LOGIC_VECTOR (3 downto 0));
    end component;
    
    component hrdata_bus_master is
         Port (
             clk : in std_logic;
             reset : in std_logic;
             hrdata_ctrl : in hrdata_ctrl_t;	
             hrdata : in std_logic_vector(31 downto 0);	
             hrdata_program_value : out std_logic_vector(31 downto 0);	
             hrdata_data_value : out std_logic_vector(31 downto 0);	
             ldm_hrdata_value : out std_logic_vector(31 downto 0);	
             SP_main_init : out std_logic_vector(31 downto 0);	
             PC_init : out std_logic_vector(31 downto 0);
             SVC_addr : out std_logic_vector(31 downto 0)	
         );
    end component;
    
    -- Declare clock interface
    ATTRIBUTE X_INTERFACE_INFO : STRING;
    ATTRIBUTE X_INTERFACE_INFO of HCLK: SIGNAL is "xilinx.com:signal:clock:1.0 HCLK CLK";
    ATTRIBUTE X_INTERFACE_PARAMETER : STRING;
    ATTRIBUTE X_INTERFACE_PARAMETER of HCLK: SIGNAL is "ASSOCIATED_RESET HRESETn, FREQ_HZ 50000000";
    
    -- Declare reset interface
    ATTRIBUTE X_INTERFACE_INFO of HRESETn: SIGNAL is "xilinx.com:signal:reset:1.0 HRESETn RST";
    ATTRIBUTE X_INTERFACE_PARAMETER of HRESETn: SIGNAL is "POLARITY ACTIVE_HIGH";

	-- M0 Core signals 
    signal PC: std_logic_vector (31 downto 0);
    signal PC_decode:  std_logic_vector (31 downto 0);
    signal PC_execute:  std_logic_vector (31 downto 0);
    signal PC_after_execute:  std_logic_vector (31 downto 0);
--	signal instruction_size : boolean;
	signal current_instruction: std_logic_vector (15 downto 0);
	signal current_instruction_32bit_HI: std_logic_vector (15 downto 0);
	signal current_instruction_final: std_logic_vector (15 downto 0);
	signal enable_decode : std_logic;
	signal data_memory_addr : std_logic_vector (31 downto 0);
	signal data_memory_addr_value : std_logic_vector (31 downto 0);
	signal hrdata_program : std_logic_vector (31 downto 0);
	signal hrdata_program_value : std_logic_vector (31 downto 0);
	signal hrdata_data : std_logic_vector (31 downto 0);
	signal hrdata_data_value : std_logic_vector (31 downto 0);
	signal hrdata_data_value_sized : std_logic_vector (31 downto 0);
	signal hrdata_data_value_16_sized : std_logic_vector (15 downto 0);
	signal ldm_hrdata_value : std_logic_vector (31 downto 0);
	signal LDM_STM_mem_address_index : unsigned (4 downto 0);
	signal LDM_STM_mem_addr : unsigned (31 downto 0);
	signal PUSH_mem_addr: unsigned (31 downto 0);
	signal POP_mem_addr: unsigned (31 downto 0);
	signal imm8_z_ext : std_logic_vector(31 downto 0) := (others => '0');			
	signal imm8_z_ext_value : std_logic_vector(31 downto 0);			
    signal internal_reset: std_logic := '1';
    signal VT_addr : std_logic_vector (31 downto 0);
	signal hrdata_NC : std_logic_vector (31 downto 0);			-- HRDATA Not Connected
	signal pos_A_is_multi_cycle : boolean;
	signal PC_plus_4 : std_logic_vector (31 downto 0);
	signal PC_after_execute_plus_4 : std_logic_vector (31 downto 0);
	signal PC_after_execute_plus_2 : std_logic_vector (31 downto 0);
	signal new_PC : std_logic_vector (31 downto 0);
	signal SDC_gp_addrB : std_logic_vector (3 downto 0);
	signal xPSR : std_logic_vector (31 downto 0);
	signal hwdara_final : std_logic_vector (31 downto 0);
	signal special_reg_content : std_logic_vector (31 downto 0);
	signal special_reg_content_value : std_logic_vector (31 downto 0);
	signal Rn : std_logic_vector (31 downto 28);
--	signal Rn_value : std_logic_vector (31 downto 28);
	signal SYSm : std_logic_vector (7 downto 0);
	signal msr_update_MSP : boolean;
	signal msr_update_PSP : boolean;
	signal msr_update_PRIMASK : boolean;
	signal msr_update_CONTROL : boolean;

	
	
   
	-- Registers after decoder
	signal gp_WR_addr : std_logic_vector(3 downto 0) := (others => '0');	
	signal gp_WR_addr_value : std_logic_vector(3 downto 0) := (others => '0');	
	signal gp_WR_addr_final : std_logic_vector(3 downto 0) := (others => '0');
    signal gp_WR_addr_non_xxM : std_logic_vector(3 downto 0) := (others => '0');	
	signal gp_addrA : std_logic_vector(3 downto 0) := (others => '0');	
	signal gp_addrB : std_logic_vector(3 downto 0) := (others => '0');			
	signal gp_addrC : std_logic_vector(3 downto 0) := (others => '0');			
	signal gp_addrA_value : std_logic_vector(3 downto 0);			
	signal gp_addrB_value : std_logic_vector(3 downto 0);			
	signal gp_addrC_value : std_logic_vector(3 downto 0);			
	signal gp_addrB_final : std_logic_vector(3 downto 0);			
	signal gp_ram_dataA : std_logic_vector(31 downto 0);			
	signal gp_ram_dataB : std_logic_vector(31 downto 0);	
	signal gp_ram_dataC : std_logic_vector(31 downto 0);	
	signal gp_addrA_executor : std_logic_vector(31 downto 0);	
	signal gp_data_in : std_logic_vector(31 downto 0);	
    signal branch_target_address : std_logic_vector (31 downto 0);
	signal branch_target_address_value : std_logic_vector (31 downto 0);
	signal prev_inst32_fields : std_logic_vector (10 downto 0);
	
   
    -- decoder signals
    signal inst32_detected_value : boolean;
    signal inst32_detected_in_prev_inst : boolean;
    signal imm8 : std_logic_vector (7 downto 0);
    signal LR_PC : std_logic;	
	signal WE : std_logic;	
	signal use_PC : boolean;
    signal access_mem : boolean;
    signal access_mem_value : boolean;
	signal PC_updated : boolean;	
	signal use_base_register : boolean;	
	signal use_base_register_value : boolean;	
	signal mem_load_size : mem_op_size_t;	
	signal mem_load_size_value : mem_op_size_t;	
	signal mem_load_sign_ext : boolean;
	signal mem_load_sign_ext_value : boolean;
	signal LDM_STM_access_mem : boolean;
	signal LDM_STM_access_mem_value : boolean;
	signal access_mem_mode : access_mem_mode_t;
	signal cond : std_logic_vector (3 downto 0);
	signal prev_inst : std_logic_vector (15 downto 0);
	
	
	-- executor signals
    signal command:  executor_cmds_t := NOT_DEF;
    signal command_value:  executor_cmds_t := NOT_DEF;
    signal result:  std_logic_vector (31 downto 0);
	signal cmd_out : executor_cmds_t;	
	signal set_flags : boolean;
	signal msr_flags : boolean;
	signal SP_updated : boolean;
	
	
	signal mem_access_exec : boolean;
	signal alu_temp_32 : std_logic;
	signal overflow_status : std_logic_vector (2 downto 0);
	signal data_mem_addr_out : std_logic_vector (31 downto 0);
	signal executor_opernd_B : std_logic_vector (31 downto 0);
	
	-- core state signals
	signal HADDR_temp  :  std_logic_vector (31 downto 0);
    signal flags       :  flag_t;
    signal instr_ptr : std_logic;
    signal disable_fetch : boolean;
    signal gp_data_in_ctrl : gp_data_in_ctrl_t;
    signal hrdata_ctrl : hrdata_ctrl_t;
    signal haddr_ctrl : haddr_ctrl_t;
    signal disable_executor : boolean;
    signal gp_addrA_executor_ctrl : boolean;
    signal LDM_W_STM_R_reg :std_logic_vector (3 downto 0);
    signal LDM_STM_capture_base : boolean;
    signal SP_main:  std_logic_vector (31 downto 0);
    signal SP_process:  std_logic_vector (31 downto 0);
    signal SP_main_init:  std_logic_vector (31 downto 0);
    signal PC_init:  std_logic_vector (31 downto 0);
    signal SVC_addr:  std_logic_vector (31 downto 0);
    signal VT_ctrl : VT_ctrl_t;
    signal SDC_push_read_address : SDC_push_read_address_t;
    signal PRIMASK:  std_logic_vector (0 downto 0);
    signal CONTROL:  std_logic_vector (1 downto 0);
    signal new_SP: std_logic_vector (31 downto 0); 
    
    
   
    signal data_memory_addr_i : unsigned (31 downto 0);
    signal LDR_mul_result : unsigned (7 downto 0);
    signal LDR_mul_result_value : unsigned (7 downto 0);
    signal LDR_multiplier : unsigned (7 downto 0);
    signal base_reg_content : std_logic_vector (31 downto 0);
    signal base_reg_content_LDM_STM : std_logic_vector (31 downto 0);
    signal mem_index_content : std_logic_vector (31 downto 0);
    signal forward_alu_result : boolean;
  
    -- pipeline_invalidator signals

    -- aliases
    -- Little endian:
    -- [      inst A 1st half    ] [     inst A 2nd half     ] [    inst B 1st half    ]   [ inst B 2nd half ] 
    -- [31 30 29 28 - 27 26 25 24] [23 22 21 20 - 19 18 17 16] [15 14 13 12 - 11 10 9 8] - [7 6 5 4 - 3 2 1 0]
    
    alias inst_A_1st_half : std_logic_vector(7 downto 0) is hrdata_program (31 downto 24);
    alias inst_A_2nd_half : std_logic_vector(7 downto 0) is hrdata_program (23 downto 16);
    alias inst_B_1st_half : std_logic_vector(7 downto 0) is hrdata_program (15 downto 8);
    alias inst_B_2nd_half : std_logic_vector(7 downto 0) is hrdata_program (7 downto 0);
    alias opcode: STD_LOGIC_VECTOR (5 downto 0) is current_instruction (15 downto 10);               -- bits (15 downto 10)
    
--    alias f32_inst_A_1st_half : std_logic_vector(7 downto 0) is fetched_32_bit_instruction (31 downto 24);
--    alias f32_inst_A_2nd_half : std_logic_vector(7 downto 0) is fetched_32_bit_instruction (23 downto 16);
--    alias f32_inst_B_1st_half : std_logic_vector(7 downto 0) is fetched_32_bit_instruction (15 downto 8);
--    alias f32_inst_B_2nd_half : std_logic_vector(7 downto 0) is fetched_32_bit_instruction (7 downto 0);
    
     signal number_of_ones_initial :  STD_LOGIC_VECTOR (3 downto 0);
     signal LDM_total_bytes_read :  STD_LOGIC_VECTOR (4 downto 0);    -- cannot exceed 7 * 4 = 28 bytes
  
	-- Simulation signals  
	--synthesis translate off
    signal cortex_m0_opcode : string(1 to 17) := "                 ";
    signal cortex_m0_status : string(1 to 18) := "NN,NZ,NC,NV, -----";
	--synthesis translate on

begin

    m0_registers: registers port map (
                            clk => HCLK,
                          reset => internal_reset,
                             WE => WE,
                     gp_WR_addr => gp_WR_addr_final, 
                     gp_data_in => gp_data_in,
                       gp_addrA => gp_addrA,
                       gp_addrB => gp_addrB_final,
                       gp_addrC => gp_addrC, 
                   gp_ram_dataA => gp_ram_dataA,
                   gp_ram_dataB => gp_ram_dataB,
                   gp_ram_dataC => gp_ram_dataC
    );
    
    m0_decoder: decoder port map ( 
                                clk => HCLK,    
                              reset => internal_reset,
                        instruction => current_instruction_final,
       inst32_detected_in_prev_inst => inst32_detected_in_prev_inst,
                    inst32_detected => inst32_detected_value,
                  destination_is_PC => PC_updated,
                         gp_WR_addr => gp_WR_addr_value,
                           gp_addrA => gp_addrA_value,
                           gp_addrB => gp_addrB_value,
                           gp_addrC => gp_addrC_value,
                               imm8 => imm8,
                              LR_PC => LR_PC,
                      execution_cmd => command_value,
                         access_mem => access_mem_value,
                  use_base_register => use_base_register_value,
                      mem_load_size => mem_load_size_value,
                  mem_load_sign_ext => mem_load_sign_ext_value,
                 LDM_STM_access_mem => LDM_STM_access_mem_value,
                    access_mem_mode => access_mem_mode,
                               cond => cond,
                          prev_inst => prev_inst
        );
    
     m0_executor: executor port map (
                            clk => HCLK,
                          reset => internal_reset,
                      operand_A => gp_addrA_executor,	
                      operand_B => executor_opernd_B,	
                        command => command, 	
                     imm8_z_ext => imm8_z_ext,
              destination_is_PC => PC_updated,
                  current_flags => flags,
                     access_mem => access_mem,
                gp_data_in_ctrl => gp_data_in_ctrl, 
               disable_executor => disable_executor,
                        SP_main => SP_main,
                        cmd_out => cmd_out,
                      set_flags => set_flags,
                         result => result,
                    alu_temp_32 => alu_temp_32,
                overflow_status => overflow_status,
                             WE => WE,
                     SP_updated => SP_updated
         );
         
      m0_core_state_m: core_state port map (
                            clk => HCLK,
                          reset => internal_reset,
--               instruction_size => instruction_size,
                     access_mem => access_mem_value,
                     PC_updated => PC_updated,
                           cond => cond,
                  current_flags => flags,
                           imm8 => imm8_z_ext(7 downto 0),
                     imm8_value => imm8_z_ext_value(7 downto 0),
              imm11_10_downto_8 => imm8_z_ext(10 downto 8),
        imm11_value_10_downto_8 => imm8_z_ext_value(10 downto 8),
                          LR_PC => LR_PC,
         number_of_ones_initial => number_of_ones_initial,
            execution_cmd_value => command_value,
             LDM_STM_access_mem => LDM_STM_access_mem_value,
                         new_PC => new_PC, 
                access_mem_mode => access_mem_mode,
                   SP_main_init => SP_main_init,
                        PC_init => PC_init,
           pos_A_is_multi_cycle => pos_A_is_multi_cycle,
               ldm_hrdata_value => ldm_hrdata_value,
          inst32_detected_value => inst32_detected_value,
   current_instruction_32bit_HI => current_instruction_32bit_HI,
            current_instruction => current_instruction_final,
                 msr_update_MSP => msr_update_MSP,
                 msr_update_PSP => msr_update_PSP,
             msr_update_PRIMASK => msr_update_PRIMASK,
             msr_update_CONTROL => msr_update_CONTROL,
                    new_PRIMASK => gp_ram_dataB (0 downto 0),
                    new_CONTROL => gp_ram_dataB (1 downto 0),
                         new_SP => new_SP,
                     SP_updated => SP_updated,
                             PC => PC,
                        SP_main => SP_main,
                     SP_process => SP_process,
                      PC_decode => PC_decode,
                     PC_execute => PC_execute,
               PC_after_execute => PC_after_execute,
      LDM_STM_mem_address_index => LDM_STM_mem_address_index,
                gp_data_in_ctrl => gp_data_in_ctrl,
                    hrdata_ctrl => hrdata_ctrl,
                  disable_fetch => disable_fetch,
                     haddr_ctrl => haddr_ctrl,
               disable_executor => disable_executor,
         gp_addrA_executor_ctrl => gp_addrA_executor_ctrl,
                LDM_W_STM_R_reg => LDM_W_STM_R_reg,
           LDM_STM_capture_base => LDM_STM_capture_base,
                         HWRITE => HWRITE,
                        VT_ctrl => VT_ctrl,
          branch_target_address => branch_target_address,
      branch_target_address_val => branch_target_address_value,
          SDC_push_read_address => SDC_push_read_address,
                inst32_detected => inst32_detected_in_prev_inst,
                             Rn => Rn,
                        PRIMASK => PRIMASK,
                        CONTROL => CONTROL
        ); 
        
     m0_core_flags: status_flags port map (
                            clk => HCLK,
                          reset => internal_reset,
                         result => result,
                           C_in => alu_temp_32,
                            cmd => cmd_out,
                      set_flags => set_flags,
                      msr_flags => msr_flags,
                     Rn_content => gp_ram_dataB (31 downto 28),
                overflow_status => overflow_status,
                       flags_o  => flags,
                           xPSR => xPSR
        );
        
     msr_flags_p : process (gp_data_in_ctrl) begin
        if (gp_data_in_ctrl = sel_Rn) and (SYSm(7 downto 3) = B"0_0000")  then
            msr_flags <= true;    
        else
            msr_flags <= false;
        end if;
     end process; 
     
     msr_update_MSP_p : process (gp_data_in_ctrl) begin
        if (gp_data_in_ctrl = sel_Rn) and (SYSm(7 downto 3) = B"0_0001" and SYSm(2 downto 0) = B"000")  then
            msr_update_MSP <= true;    
        else
            msr_update_MSP <= false;
        end if;
     end process;  
     
      msr_update_PSP_p : process (gp_data_in_ctrl) begin
        if (gp_data_in_ctrl = sel_Rn) and (SYSm(7 downto 3) = B"0_0001" and SYSm(2 downto 0) = B"001")  then
            msr_update_PSP <= true;    
        else
            msr_update_PSP <= false;
        end if;
     end process;  
     
     msr_update_PRIMASK_p : process (gp_data_in_ctrl) begin
        if (gp_data_in_ctrl = sel_Rn) and (SYSm(7 downto 3) = B"0_0010" and SYSm(2 downto 0) = B"000")  then
            msr_update_PRIMASK <= true;    
        else
            msr_update_PRIMASK <= false;
        end if;
     end process;  
     
     msr_update_CONTROL_p : process (gp_data_in_ctrl) begin
        if (gp_data_in_ctrl = sel_Rn) and (SYSm(7 downto 3) = B"0_0010" and SYSm(2 downto 0) = B"100")  then
            msr_update_CONTROL <= true;    
        else
            msr_update_CONTROL <= false;
        end if;
     end process;  
        
     m0_count_ones: count_ones port map ( 
                        byte_in => imm8_z_ext(7 downto 0),
                           ones => number_of_ones_initial
        );    
        
     hrdata_bus_master_m0: hrdata_bus_master  port map (
             clk => HCLK,
             reset => internal_reset,
             hrdata_ctrl => hrdata_ctrl,
             hrdata => HRDATA, 
             hrdata_program_value => hrdata_program_value,
             hrdata_data_value => hrdata_data_value,
             ldm_hrdata_value => ldm_hrdata_value,
             SP_main_init => SP_main_init,
             PC_init => PC_init,
             SVC_addr => SVC_addr
         );
        
    LDM_total_bytes_read <= std_logic_vector (shift_left(unsigned('0' & number_of_ones_initial), 2)); --   
    PC_plus_4 <= std_logic_vector ((unsigned (PC) + 4));
    
    new_PC_p : process (result, command, gp_ram_dataA, SVC_addr, haddr_ctrl) begin
        if (haddr_ctrl = sel_SVC_mem_content) then
            new_PC <= SVC_addr; 
        elsif (command = BX or command = BLX) then
            new_PC <= gp_ram_dataA;   
        else
            new_PC <= result;
        end if;
    end process;
    
    new_SP_p : process (gp_ram_dataB, result, SP_updated) begin
        if (SP_updated) then
            new_SP <= result; 
        else
            new_SP <= gp_ram_dataB; 
        end if;
    end process;
  
    pos_A_is_multi_cycle_p : process (HCLK, internal_reset) begin
       if (internal_reset = '1') then
           pos_A_is_multi_cycle <= false;
       else
           if (rising_edge (HCLK)) then
                if (PC(1) = '0') then
                    -- instruction at position A
                    if (command_value = LDR_imm5 or 
                        command_value = LDR_SP_imm8 or 
                        command_value = LDRH_imm5 or 
                        command_value = LDRB_imm5 or 
                        command_value = LDR or 
                        command_value = LDRH or 
                        command_value = LDRSH or 
                        command_value = LDRB or 
                        command_value = LDRSB or 
                        command_value = LDM or 
                        command_value = STR_imm5 or 
                        command_value = STRH_imm5 or 
                        command_value = STRB_imm5 or 
                        command_value = STR or 
                        command_value = STRH or 
                        command_value = STRB or 
                        command_value = STR_SP_imm8 or 
                        command_value = STM or 
                        command_value = PUSH or 
                        command_value = POP or
                        command_value = EVAL_32_INSTR   
                        ) then
                        pos_A_is_multi_cycle <= true;
                    else
                        pos_A_is_multi_cycle <= false;    
                    end if;
                end if;      
           end if;                       
       end if;
    end process;  
        
    ---------------------------------------------------------------------------------------
    --- Hardware which drives (Cortex-M0) module input/ouput pins
    ---------------------------------------------------------------------------------------    
    
    HWDATA <= hwdara_final;
    
    HSIZE_p : process (mem_load_size) begin
        case (mem_load_size) is
            when WORD           =>  HSIZE <= "010";
            when HALF_WORD      =>  HSIZE <= "001";  
            when BYTE           =>  HSIZE <= "000";  
            when others         =>  null;  
        end case; 
    end process;  
    
    VT_addr_p : process (VT_ctrl) begin
        case (VT_ctrl) is                                           -- Vector Table index
            when    VT_SP_main =>  VT_addr <= x"0000_0000";         -- 0
            when      VT_RESET =>  VT_addr <= x"0000_0004";         -- 1
            when        VT_NMI =>  VT_addr <= x"0000_0008";         -- 2
            when  VT_HardFault =>  VT_addr <= x"0000_000C";         -- 3
            when     VT_SVCall =>  VT_addr <= x"0000_002C";         -- 11
            when     VT_PendSV =>  VT_addr <= x"0000_0038";         -- 14
            when    VT_SysTick =>  VT_addr <= x"0000_003C";         -- 15
            when       VT_NONE =>  VT_addr <= x"0000_0000";
            when others        =>   null;  
        end case; 
    end process;  
      
    hwdara_final_p : process (SDC_push_read_address, PC_execute, xPSR, gp_ram_dataB) begin
         case (SDC_push_read_address) is
            when SDC_read_retuen_addr     => hwdara_final <= PC_execute;
            when SDC_read_xPSR            => hwdara_final <= xPSR;
            when others                   => hwdara_final <= gp_ram_dataB;
        end case;
    end process;     
  
    
    HADDR_temp_p : process ( LDM_STM_access_mem, haddr_ctrl, data_memory_addr, data_memory_addr_i, 
                        PC(31 downto 2), LDM_STM_mem_addr, VT_addr, PUSH_mem_addr, POP_mem_addr, 
                        branch_target_address_value, branch_target_address, new_PC, SVC_addr) begin
--        if (command_value = SVC) then        
--            HADDR <= x"0000_002C";      -- SVC exception no. = 11 * 4 = 44 = 0x2C 
--        else                
            case (haddr_ctrl) is
                when              sel_PC         =>  HADDR_temp <= PC(31 downto 2) & B"00";  
                when            sel_DATA         =>  HADDR_temp <= data_memory_addr;
                when             sel_LDM         =>  HADDR_temp <= std_logic_vector (LDM_STM_mem_addr);
                when             sel_STM         =>  HADDR_temp <= std_logic_vector (LDM_STM_mem_addr);
                when           sel_WDATA         =>  HADDR_temp <= std_logic_vector (data_memory_addr_i);
                when    sel_VECTOR_TABLE         =>  HADDR_temp <= VT_addr;
                when    sel_SP_main_addr         =>  HADDR_temp <= std_logic_vector (PUSH_mem_addr);
                when    sel_SP_main_addr_plus_4  =>  HADDR_temp <= std_logic_vector (POP_mem_addr);
                when       sel_PC_plus_4         =>  HADDR_temp <=  PC_plus_4 (31 downto 2) & B"00";  
                when          sel_BRANCH         =>  HADDR_temp <= std_logic_vector (branch_target_address_value);
                when       sel_BRANCH_BL         =>  HADDR_temp <= std_logic_vector (branch_target_address);
                when           sel_BX_Rm         =>  HADDR_temp <= new_PC;
                when          sel_BLX_Rm         =>  HADDR_temp <= new_PC;
                when    sel_SP_main_addr_SVC     =>  HADDR_temp <= std_logic_vector (PUSH_mem_addr);
                when    sel_SVC_mem_content      =>  HADDR_temp <= SVC_addr;
                when        others               =>  null;
            end case;
--        end if;
    end process;   
    
    HADDR <= HADDR_temp;
   
    LDM_STM_mem_addr <= (unsigned (base_reg_content_LDM_STM) + LDM_STM_mem_address_index) and x"FFFF_FFFE";     -- gp_ram_dataA holds the base value (Rn)
    PUSH_mem_addr <=  unsigned (SP_main and x"FFFF_FFFE");
    POP_mem_addr <=   unsigned ((unsigned (SP_main) + 4) and x"FFFF_FFFE");
    
  
    internal_reset <= not HRESETn;
    HBURST <= B"000";
    HMASTLOCK <= '0';
    HPROT <= B"0000";
    HPROT <= B"0000";
    HTRANS <= B"00";
    
    ---------------------------------------------------------------------------------------
    --- Hardware which drives (Executor) module input pins
    ---------------------------------------------------------------------------------------
    
    gp_addrA_executor_p: process (gp_ram_dataA, hrdata_data, access_mem, 
                                  gp_addrA_executor_ctrl, PC_after_execute) begin
        if (access_mem = true) then       -- Desitinatination register is PC
            gp_addrA_executor <= hrdata_data;        
        else
            if (gp_addrA_executor_ctrl = true) then       -- Desitinatination register is PC
                gp_addrA_executor <= PC_after_execute;        
            else
                gp_addrA_executor <= gp_ram_dataA;
            end if;
        end if;        
    end process;

    executor_opernd_B_p: process (gp_ram_dataB, access_mem, PC) begin
        if (access_mem = true) then
             executor_opernd_B <= PC;  
        else
             executor_opernd_B <= gp_ram_dataB;
        end if;   
    end process; 
    
    ---------------------------------------------------------------------------------------
    --- Hardware which drives (Register) module input pins
    ---------------------------------------------------------------------------------------
    
    special_reg_content_value_p : process (imm8, flags, SP_main) begin
        case (imm8) is
            when sp_reg_APSR =>  special_reg_content_value <=                -- The flags from previous instructions.
                to_std_logic (flags.N) &        -- bit 31
                to_std_logic (flags.Z) &        -- bit 30
                to_std_logic (flags.C) &        -- bit 29
                to_std_logic (flags.V) &        -- bit 28
                x"0_00_0000";        
            when sp_reg_IAPSR =>  special_reg_content_value <=                -- A composite of IPSR and APSR.
                to_std_logic (flags.N) &        -- bit 31
                to_std_logic (flags.Z) &        -- bit 30
                to_std_logic (flags.C) &        -- bit 29
                to_std_logic (flags.V) &        -- bit 28
                x"0_00_00" & B"00" &
                to_std_logic_vector (flags.EN); -- bit 5 downto 0   
            when sp_reg_EAPSR =>  special_reg_content_value <=                -- A composite of EPSR and APSR.
                to_std_logic (flags.N) &        -- bit 31
                to_std_logic (flags.Z) &        -- bit 30
                to_std_logic (flags.C) &        -- bit 29
                to_std_logic (flags.V) &        -- bit 28
                B"000" &
                to_std_logic (flags.T) &        -- bit 24
                x"00_0000";
            when sp_reg_XPSR =>  special_reg_content_value <=                 -- A composite of all three PSR registers.
                to_std_logic (flags.N) &        -- bit 31
                to_std_logic (flags.Z) &        -- bit 30
                to_std_logic (flags.C) &        -- bit 29
                to_std_logic (flags.V) &        -- bit 28   
                B"000" &
                to_std_logic (flags.T) &        -- bit 24   
                x"0000" & B"00" &
                to_std_logic_vector (flags.EN); -- bit 5 downto 0   
            when sp_reg_IPSR =>  special_reg_content_value <=                 -- The Interrupt status register.
                x"00_0000" & B"00" &
                to_std_logic_vector (flags.EN); -- bit 5 downto 0   
            when sp_reg_EPSR =>  special_reg_content_value <=                 -- The execution status register.
                x"0" &
                B"000" &
                to_std_logic (flags.T) &        -- bit 24
                x"00_0000";
            when sp_reg_IEPSR =>  special_reg_content_value <=                 -- A composite of IPSR and EPSR.
                x"0" &
                B"000" &
                to_std_logic (flags.T) &        -- bit 24
                x"0000" & B"00" &
                to_std_logic_vector (flags.EN); -- bit 5 downto 0   
            when sp_reg_MSP =>  special_reg_content_value <=                   -- The Main Stack pointer.
                SP_main;    
            when sp_reg_PSP =>  special_reg_content_value <=                   -- The Process Stack pointer.
                SP_main;                        -- TODO: Process Stack pointer not yet implemented.
            when sp_reg_PRIMASK =>  special_reg_content_value <=               -- Register to mask out configurable exceptions.
                x"0000000" & B"000" &
                PRIMASK; 
            when sp_reg_CONTROL =>  special_reg_content_value <=               -- The CONTROL register.
                 x"000_0000" & B"00" &
                 CONTROL;
            when others =>  special_reg_content_value <=
                x"0000_0000";                                                                         
        end case; 
    end process;
    
    SDC_gp_addrB_p : process (SDC_push_read_address) begin
        case (SDC_push_read_address) is
            when SDC_read_R0            => SDC_gp_addrB <= B"0000";
            when SDC_read_R1            => SDC_gp_addrB <= B"0001";
            when SDC_read_R2            => SDC_gp_addrB <= B"0010";
            when SDC_read_R3            => SDC_gp_addrB <= B"0011";
            when SDC_read_R12           => SDC_gp_addrB <= B"1100";
            when SDC_read_R14           => SDC_gp_addrB <= B"1110";
            when SDC_read_retuen_addr   => SDC_gp_addrB <= B"0000";
            when SDC_read_xPSR          => SDC_gp_addrB <= B"0000";
            when others                 => SDC_gp_addrB <= B"0000";
        end case;
    end process;
    
    gp_WR_addr_non_xxM_p: process (haddr_ctrl, gp_WR_addr) begin
        if (haddr_ctrl = sel_BLX_Rm) then
            gp_WR_addr_non_xxM <= B"1110";           -- LR register
        else
            gp_WR_addr_non_xxM <= gp_WR_addr;
        end if;    
    end process;
    
     gp_WR_addr_final_p: process (LDM_STM_access_mem, LDM_W_STM_R_reg, disable_executor, gp_AddrA, gp_WR_addr_non_xxM) begin
         if (LDM_STM_access_mem = true) then
            if (disable_executor = true) then 
                gp_WR_addr_final <= gp_AddrA;       -- Save the Rn in LDM instruction into gp_AddrA register.
            else 
                gp_WR_addr_final <= LDM_W_STM_R_reg;
            end if;  
         else
            gp_WR_addr_final <= gp_WR_addr_non_xxM;
         end if;   
    end process;
    
    PC_after_execute_plus_4 <= std_logic_vector (unsigned (PC_after_execute) + 4);
    PC_after_execute_plus_2 <= std_logic_vector (unsigned (PC_after_execute) + 2);    
    
    gp_data_in_p: process (gp_data_in_ctrl, result, hrdata_data_value_sized, ldm_hrdata_value, 
                            PC_after_execute, LDM_total_bytes_read, gp_ram_dataA, special_reg_content) begin
        case (gp_data_in_ctrl) is 
            when sel_ALU_RESULT             => gp_data_in <= result;
            when sel_HRDATA_VALUE_SIZED     => gp_data_in <= hrdata_data_value_sized;  
            when sel_LDM_DATA               => gp_data_in <= ldm_hrdata_value;
            when sel_LDM_Rn                 => gp_data_in <= std_logic_vector (unsigned (gp_ram_dataA) + unsigned (LDM_total_bytes_read));
            when sel_SP_main_init           => gp_data_in <= result;
            when sel_PC_init                => gp_data_in <= result;
            when sel_STM_total_bytes_wrote  => gp_data_in <= std_logic_vector (unsigned (gp_ram_dataA) + unsigned (LDM_total_bytes_read));
            when sel_gp_data_in_NC          => gp_data_in <= (others => '0');
            when sel_SP_set                 => gp_data_in <= (others => '0');
            when sel_LR_DATA_BL             => gp_data_in <= PC_after_execute_plus_2(31 downto 1) & '1';
            when sel_LR_DATA_BLX            => gp_data_in <= PC_after_execute_plus_2(31 downto 1) & '1';
            when sel_special_reg            => gp_data_in <= special_reg_content;
            when sel_Rn                     => gp_data_in <= (others => '0');
            when others                     => gp_data_in <= (others => '0'); report " gp_data_in error" severity failure;
        end case;
    end process;
    
    gp_addrB_final_p: process (haddr_ctrl, use_base_register, gp_addrB_value, gp_addrB, 
                                LDM_W_STM_R_reg, SDC_gp_addrB, msr_flags, Rn, msr_update_MSP,
                                msr_update_PSP, msr_update_PRIMASK, msr_update_CONTROL) begin
        if msr_flags or msr_update_MSP or msr_update_PSP or msr_update_PRIMASK or msr_update_CONTROL  then
            gp_addrB_final <= Rn;         
        else                   
            if (haddr_ctrl = sel_STM or haddr_ctrl = sel_SP_main_addr) then
                gp_addrB_final <= LDM_W_STM_R_reg;   
            elsif (haddr_ctrl = sel_SP_main_addr_SVC) then    
                gp_addrB_final <= SDC_gp_addrB; 
            else
                if (use_base_register = true) then 
                     gp_addrB_final <= gp_addrB_value;  
                else
                     gp_addrB_final <= gp_addrB;
                end if;
            end if;   
        end if;  
    end process;
    
    
    hrdata_data_value_sized_p: process (mem_load_size, mem_load_sign_ext, hrdata_data_value, 
                                        hrdata_data_value_16_sized, data_memory_addr_i(1 downto 0)) 
        variable case_sel: unsigned (1 downto 0);
    begin
        case_sel := data_memory_addr_i (1 downto 0);
        case (mem_load_size) is
            when WORD       => hrdata_data_value_sized <= hrdata_data_value;
            when HALF_WORD  => 
                if (mem_load_sign_ext = true) then
                    if (hrdata_data_value_16_sized(15) = '1') then
                        -- negative sign extension
                        hrdata_data_value_sized <= x"FFFF" & hrdata_data_value_16_sized;    
                    else
                        hrdata_data_value_sized <= x"0000" & hrdata_data_value_16_sized;
                    end if;        
                else
                    hrdata_data_value_sized <= x"0000" & hrdata_data_value_16_sized;
                end if;
            when BYTE       =>
                if (mem_load_sign_ext = true) then
                    case (case_sel) is
                        when B"00" => hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (7 downto 0);
                        when B"01" => hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (15 downto 8);
                        when B"10" => hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (23 downto 16);
                        when B"11" => hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (31 downto 24);
                        when others =>
                            null;
                    end case;   
                else
                    case (case_sel) is
                        when B"00" => 
                            if (hrdata_data_value(7) = '0') then 
                                hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (7 downto 0);
                            else
                                hrdata_data_value_sized <=  x"FFFF_FF" & hrdata_data_value (7 downto 0);
                            end if;
                        when B"01" =>
                            if (hrdata_data_value(15) = '0') then 
                                hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (15 downto 8);
                            else
                                hrdata_data_value_sized <=  x"FFFF_FF" & hrdata_data_value (15 downto 8);
                            end if;
                        when B"10" => 
                            if (hrdata_data_value(23) = '0') then 
                                hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (23 downto 16);
                            else
                                hrdata_data_value_sized <=  x"FFFF_FF" & hrdata_data_value (23 downto 16);
                            end if;   
                        when B"11" => 
                            if (hrdata_data_value(31) = '0') then 
                                hrdata_data_value_sized <=  x"0000_00" & hrdata_data_value (31 downto 24);
                            else
                                hrdata_data_value_sized <=  x"FFFF_FF" & hrdata_data_value (31 downto 24);
                            end if;   
                        when others =>
                            null;
                    end case;  
                end if;
            when NOT_DEF    => hrdata_data_value_sized <= hrdata_data_value;
        end case;
    end process;

    hrdata_data_value_16_sized_p: process (hrdata_data_value, data_memory_addr_i(1)) begin
        if (data_memory_addr_i(1) = '1') then
            hrdata_data_value_16_sized <= hrdata_data_value (31 downto 16);      -- High Half Word
        else
            hrdata_data_value_16_sized <= hrdata_data_value (15 downto 0);       -- Low Half Word
        end if;    
    end process;
    
   
   

    
    ---------------------------------------------------------------------------------------
    --- Hardware which drives (Decoder)
    ---------------------------------------------------------------------------------------     
    current_instruction_p: process (PC(1), hrdata_program) begin
        if (PC(1) = '0') then
            current_instruction <= hrdata_program(31 downto 16);    
        else    
            current_instruction <= hrdata_program(15 downto 0);    
        end if;
    end process;
    
  
    flipflops_32bit_instruction_p: process (HCLK, internal_reset) begin
        if (internal_reset = '1') then
            current_instruction_32bit_HI <= (others => '0');
        else
            if (rising_edge (HCLK)) then
  
                if (command_value = EVAL_32_INSTR) then
                    current_instruction_32bit_HI <= current_instruction;
                end if;    
            end if;
        end if;
    end process;
    
--    current_instruction_final_p: process (is_32bit_instruction, current_instruction_32bit_HI, current_instruction) begin
--        if (is_32bit_instruction = true) then
--            current_instruction_final <= current_instruction_32bit_HI;
--        else
--            current_instruction_final <= current_instruction;
--        end if;       
--    end process;

    current_instruction_final <= current_instruction;

    imm8_z_ext_value_p: process  (command_value, gp_addrA_value, imm8) begin
        case (command_value) is
            when MOVS_imm8      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when ADDS_imm3      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when ADDS_imm8      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when ADD_SP_imm8    => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when SUBS_imm3      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when SUBS_imm8      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when SUB_SP_imm7    => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when CMP_imm8       => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LSLS_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LSRS_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when ASRS_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LDR_imm5       => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LDR_SP_imm8    => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LDRH_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LDRB_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LDR_label      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when LDM            => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when STR_imm5       => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when STRH_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when STRB_imm5      => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when STR_SP_imm8    => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when STM            => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when PUSH           => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when POP            => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when BRANCH         => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when BRANCH_imm11   => imm8_z_ext_value <= x"0000_0" & '0' & gp_addrA_value(2 downto 0) & imm8;  -- Zero extend
            when BL             => imm8_z_ext_value <= x"0000_0" & '0' & gp_addrA_value(2 downto 0) & imm8;  -- Zero extend
            when CPS            => imm8_z_ext_value <= x"0000_00" & imm8;  -- Zero extend
            when ADD_SP_SP_imm7 => imm8_z_ext_value <= x"0000_0" & B"00" & imm8 & B"00";  -- Zero extend
            when others  => imm8_z_ext_value <= (others => '0');
        end case;       
    end process; 
    
    -- data_memory_addr_value
    ----------------------------------------------------------------------------------------  
    LDR_multiplier_p: process (mem_load_size_value) begin
         case (mem_load_size_value) is
            when WORD       => LDR_multiplier <= x"02";
            when HALF_WORD  => LDR_multiplier <= x"01";
            when BYTE       => LDR_multiplier <= x"00";
            when NOT_DEF    => LDR_multiplier <= x"02";
        end case;
    end process;
    
    LDR_mul_result_value_p: process (command_value, imm8, LDR_multiplier, mem_index_content(7 downto 0), 
                                     PC_execute, LDR_mul_result_value) 
        --variable calc_index : unsigned (7 downto 0);        -- Calculate index by dividing : Word: divide by 4, HWord: divide by 2, Byte: no change                             
                                     begin
        case (command_value) is
            when LDR_imm5 | LDR_SP_imm8 | LDRH_imm5 | LDRB_imm5 | LDR_label | STR_imm5 | STRH_imm5 | STRB_imm5 | STR_SP_imm8  => 
                LDR_mul_result_value <= shift_left (unsigned (imm8), to_integer(LDR_multiplier));
            when LDR | LDRH | LDRSH | LDRB | LDRSB =>
                LDR_mul_result_value <= shift_left (unsigned (mem_index_content(7 downto 0)), to_integer(LDR_multiplier));     
            when STR =>
                --calc_index := shift_right (unsigned (mem_index_content(7 downto 0)), 2); -- Divide by 4
                --LDR_mul_result_value <= shift_left (calc_index, to_integer(LDR_multiplier));  
                LDR_mul_result_value <=  unsigned (mem_index_content(7 downto 0));  
            when STRH =>
                --calc_index := shift_right (unsigned (mem_index_content(7 downto 0)), 1); -- Divide by 2
                --LDR_mul_result_value <= shift_left (calc_index, to_integer(LDR_multiplier));    
                LDR_mul_result_value <=  unsigned (mem_index_content(7 downto 0));  
            when STRB =>
                -- No change
                --LDR_mul_result_value <= shift_left (unsigned (mem_index_content(7 downto 0)), to_integer(LDR_multiplier));   
                LDR_mul_result_value <=  unsigned (mem_index_content(7 downto 0));  

            when others =>
                null;    
        end case;
    end process; 
    
    
    forward_alu_result_p: process (gp_WR_addr, gp_addrB_final, gp_addrA_value) begin
        if (gp_WR_addr = gp_addrB_final or gp_WR_addr = gp_addrA_value) then 
            forward_alu_result <= true;
        else
            forward_alu_result <= false;
        end if;   
    end process;
    
    base_reg_content_p: process (forward_alu_result, gp_data_in, gp_ram_dataB, 
                                 gp_ram_dataA, gp_ram_dataC, gp_addrA_value, command_value, SP_main) begin
        if (forward_alu_result = true) then 
            if (gp_WR_addr = gp_addrA_value) then
                if (command_value = STR or command_value = STRH or command_value = STRB) then
                    mem_index_content <= gp_ram_dataC; 
                else
                    mem_index_content <= gp_ram_dataB; 
                end if;
                 if (command_value = STR_SP_imm8) then
                    base_reg_content <= SP_main;
                else
                   base_reg_content <= gp_data_in;  
                end if;         
            else
                if (command_value = STR or command_value = STRH or command_value = STRB) then
                    mem_index_content <= gp_ram_dataC;
                else
                    mem_index_content <= gp_data_in;
                end if;
                if (command_value = STR_SP_imm8) then
                    base_reg_content <= SP_main;
                else
                    base_reg_content <= gp_ram_dataA;  
                end if; 
            end if;    
        else
            if (command_value = STR or command_value = STRH or command_value = STRB) then
                mem_index_content <= gp_ram_dataC;
            else
                mem_index_content <= gp_ram_dataB;
            end if;
            if (command_value = STR_SP_imm8) then
                base_reg_content <= SP_main;
            else
                base_reg_content <= gp_ram_dataA;
            end if;    
            
        end if;   
    end process;
    
    base_reg_content_LDM_STM_STM_p: process (LDM_STM_capture_base, gp_ram_dataA) begin
        if (LDM_STM_capture_base = true) then
            base_reg_content_LDM_STM <= gp_ram_dataA;
        end if;   
    end process;
    
    -- TODO check to see if inserting a flip flip before use_base_register and adding use_base_register_value 
    --      breaks LDM and STM or not. 
    data_memory_addr_value_p: process (command_value, gp_ram_dataA, PC_execute, base_reg_content, 
                                       LDR_mul_result_value, use_base_register) begin
        if (use_base_register = true) then 
            if (command_value = LDM or command_value = STM) then
                data_memory_addr_i <=  unsigned (base_reg_content); -- Expected to be aligned or HardFaault
            else
                data_memory_addr_i <= unsigned (base_reg_content) +  unsigned(x"0000_00" & LDR_mul_result_value); 
            end if;    
        else
            case (command_value) is
                when LDR_label => 
                    data_memory_addr_i <= unsigned (PC_execute and x"FFFF_FFFC") +  
                                          unsigned(x"0000_00" & LDR_mul_result_value) + x"0000_0004"; 
                when LDR| LDRH | LDRSH | LDRB | STR | STRH |STRB =>
                    data_memory_addr_i <= unsigned (gp_ram_dataA) +  unsigned(x"0000_00" & LDR_mul_result_value);     
                when others =>
                        null;     
            end case;
             
        end if;   
    end process;
    
    data_memory_addr_value <= std_logic_vector (data_memory_addr_i);   
    -----------------------------------------------------------------------------------------

    decoder_registers_p: process (HCLK, internal_reset) begin 
        if internal_reset = '1' then
            imm8_z_ext <= (others => '0');
            gp_WR_addr <= (others => '0');
            gp_addrA <= (others => '0');
            gp_addrB <= (others => '0');
            gp_addrC <= (others => '0');
            command <= NOP;    
            access_mem <= false;
            hrdata_data <= (others => '0');
            hrdata_program <= (others => '0');
            data_memory_addr <= (others => '0');
            LDR_mul_result <= (others => '0');
            mem_load_sign_ext <= false;
            LDM_STM_access_mem <= false;
            use_base_register <= false;
            special_reg_content <= (others => '0');
            SYSm <= B"0000_0000";
        else
            if (rising_edge(HCLK)) then
                    imm8_z_ext <= imm8_z_ext_value;
                    gp_WR_addr <= gp_WR_addr_value;
                    gp_addrA <= gp_addrA_value;
                    gp_addrB <= gp_addrB_value;
                    gp_addrC <= gp_addrC_value;
                    command <= command_value;
                    mem_load_size <= mem_load_size_value;
                    data_memory_addr <= data_memory_addr_value;
                    LDR_mul_result <= LDR_mul_result_value;
                    mem_load_sign_ext <= mem_load_sign_ext_value;
                    LDM_STM_access_mem <= LDM_STM_access_mem_value;
                    use_base_register <= use_base_register_value;
                    special_reg_content <= special_reg_content_value;
                    SYSm <= current_instruction_final (7 downto 0);
                    if (disable_fetch = false) then
                        access_mem <= access_mem_value;
                        hrdata_data <= hrdata_data_value; 
                        hrdata_program <= hrdata_program_value;
                    end if;  
            end if;    
        end if;
    end process;
    
    
    -----------------------------------------------------------------------------------------
    -- Reconfigurable related codes start from here.
    -----------------------------------------------------------------------------------------
    
--    m0_RC_PC_sensivity_i: m0_RC_PC_sensivity port map( 
--            HADDR => HADDR_temp,
--            invoke_accelerator => invoke_accelerator
--        );


    -----------------------------------------------------------------------------------------
    -- Simulation related code starts here,
    -- These section will not be synthesized.
    -----------------------------------------------------------------------------------------
    --synthesis translate off
    
    simulation_status_p: process (HCLK, internal_reset, flags) 
    begin
      
        if rising_edge(HCLK) then 
            if internal_reset = '1' then
                cortex_m0_status <= "NN,NZ,NC,NV, Reset"; 
            else
                if (flags.N = '1') then cortex_m0_status(1 to 3)   <= " N,"; else cortex_m0_status(1 to 3)   <= "NN,"; end if;
                if (flags.Z = '1') then cortex_m0_status(4 to 6)   <= " Z,"; else cortex_m0_status(4 to 6)   <= "NZ,"; end if;
                if (flags.C = '1') then cortex_m0_status(7 to 9)   <= " C,"; else cortex_m0_status(7 to 9)   <= "NC,"; end if;
                if (flags.V = '1') then cortex_m0_status(10 to 12) <= " V,"; else cortex_m0_status(10 to 12) <= "NV,"; end if;
                cortex_m0_status(13 to 18) <= " ,Run ";
            end if;      
        end if;      
    end process;

    simulation_p: process (internal_reset, inst32_detected_in_prev_inst, inst32_detected_value, current_instruction_final, prev_inst)
        -- Variables for contents of each register in each bank
        -- variable sim_r0 : std_logic_vector(31 downto 0) := X"0000";
        variable     Rd_decode : string(1 to 2);   -- Rd register specification
        variable     Rm_decode : string(1 to 2);   -- Rd register specification
        variable     Rn_decode : string(1 to 2);   -- Rn register specification
        variable     imm8_decode : string(1 to 3);   -- immediate 8 specification
        variable     imm11_decode : string(1 to 4);   -- immediate 8 specification
        variable     LR_PC_decode : string(1 to 2);
        variable     cond_decode : string(1 to 2);
    begin  
        Rd_decode (1) := 'r';
        Rm_decode (1) := 'r';
        Rn_decode (1) := 'r';
        imm8_decode (1) :=  '#';
        imm11_decode (1) :=  '#';
        LR_PC_decode (1) := '#';
        
    if internal_reset = '1' then
        cortex_m0_opcode <= "CORE IS RESET!   ";
    else            
        if (inst32_detected_in_prev_inst = true) then
            if std_match(current_instruction_final(14 downto 12), "1-1") then
                -- BL
                imm11_decode (2) :=  hexcharacter ('0' & current_instruction_final (10 downto 8));
                imm11_decode (3) :=  hexcharacter (current_instruction_final (7 downto 4));
                imm11_decode (4) :=  hexcharacter (current_instruction_final (3 downto 0));  
                cortex_m0_opcode <= "BL" & " ,{" & imm11_decode & "}"  & "       ";  
            elsif  std_match(prev_inst(10 downto 4), "011100-") then
                -- MSR
                Rn_decode(2) := hexcharacter (prev_inst (3 downto 0));
                imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                cortex_m0_opcode <= "MSR <" & imm8_decode & ">, <" & Rn_decode & ">  ";  
            elsif  std_match(prev_inst(10 downto 4), "011111-") then
                -- MRS
                Rd_decode(2) := hexcharacter (current_instruction_final (11 downto 8));
                imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                cortex_m0_opcode <= "MRS <" & Rn_decode & ">, <" & imm8_decode & ">  ";  
            elsif  std_match(prev_inst(10 downto 4), "0111011") and std_match(current_instruction_final(7 downto 4), "0100") then
                -- DSB
                imm8_decode(2) :=  hexcharacter ("0000");
                imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                cortex_m0_opcode <= "DSB #" & imm8_decode & "         ";
            elsif  std_match(prev_inst(10 downto 4), "0111011") and std_match(current_instruction_final(7 downto 4), "0101") then
                -- DMB
                imm8_decode(2) :=  hexcharacter ("0000");
                imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                cortex_m0_opcode <= "DMB #" & imm8_decode & "         ";
            elsif  std_match(prev_inst(10 downto 4), "0111011") and std_match(current_instruction_final(7 downto 4), "0110") then
                -- ISB
                imm8_decode(2) :=  hexcharacter ("0000");
                imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                cortex_m0_opcode <= "ISB #" & imm8_decode & "         ";
            else
                -- UNKNOWN 32-bit instruction
            end if;
        else
            if (inst32_detected_value = false) then
                -------------------------------------------------------------------------------------- -- MOVS Rd, #(imm8)
                if std_match(current_instruction_final(15 downto 10), "00100-") then                      
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8));               
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "MOVS " & Rd_decode & "," & imm8_decode & "      ";    
                -------------------------------------------------------------------------------------- -- MOVS <Rd>,<Rm>     
                elsif std_match(current_instruction_final(15 downto 6), "0000000000") then                 
                    Rd_decode(2) := hexcharacter (current_instruction_final (3 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "MOVS " & Rd_decode & "," & Rm_decode & "       "; 
                -------------------------------------------------------------------------------------- -- MOV <Rd>,<Rm>  ,  MOV PC, Rm     
                elsif std_match(current_instruction_final(15 downto 8), "01000110") then                   
                    Rd_decode(2) := hexcharacter (current_instruction_final (7) & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter (current_instruction_final (6 downto 3));
                    cortex_m0_opcode <= "MOV  " & Rd_decode & "," & Rm_decode & "       ";    
                -------------------------------------------------------------------------------------- -- ADDS <Rd>,<Rn>,#<imm3>
                elsif std_match(current_instruction_final(15 downto 9), "0001110") then                    
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    imm8_decode(3) :=   hexcharacter ('0' & current_instruction_final (8 downto 6));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "ADDS " & Rd_decode & "," & Rn_decode & "," & imm8_decode & "   ";    
                -------------------------------------------------------------------------------------- -- ADDS <Rd>,<Rn>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 9), "0001100") then                   
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6));
                    cortex_m0_opcode <= "ADDS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";    
                -------------------------------------------------------------------------------------- -- ADD <Rdn>,<Rm> - ADD PC,<Rm>
                elsif std_match(current_instruction_final(15 downto 8), "01000100") then                  
                    Rd_decode(2) := hexcharacter (current_instruction_final(7) & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter (current_instruction_final (6 downto 3));
                    cortex_m0_opcode <= "ADD  " & Rd_decode & "," & Rm_decode & "       ";    
                -------------------------------------------------------------------------------------- -- ADDS <Rdn>,#<imm8>
                elsif std_match(current_instruction_final(15 downto 11), "00110") then                      
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8));
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "ADDS " & Rd_decode & "," & imm8_decode & "      ";    
                -------------------------------------------------------------------------------------- -- ADCS <Rdn>,<Rm>  
                elsif std_match(current_instruction_final(15 downto 6), "0100000101") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "ADCS " & Rd_decode & "," & Rm_decode & "       "; 
                -------------------------------------------------------------------------------------- -- ADD <Rd>,SP,#<imm8>  
                elsif std_match(current_instruction_final(15 downto 11), "10101") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8));
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "ADD " & Rd_decode & ",SP," & imm8_decode & "    ";     
                -------------------------------------------------------------------------------------- -- ADD SP,SP,#<imm8>  
                elsif std_match(current_instruction_final(15 downto 7), "101100000") then                
                    imm8_decode(2) :=   hexcharacter ('0' & current_instruction_final (6 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "ADD " & "SP,SP," & imm8_decode & "    ";
                -------------------------------------------------------------------------------------- -- SUBS <Rd>,<Rn>,#<imm3>  
                elsif std_match(current_instruction_final(15 downto 9), "0001111") then                  
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    imm8_decode(3) :=   hexcharacter ('0' & current_instruction_final (8 downto 6));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "SUBS " & Rd_decode & "," & Rn_decode & "," & imm8_decode & "   ";  
                -------------------------------------------------------------------------------------- -- SUBS <Rd>,<Rn>,<Rm>  
                elsif std_match(current_instruction_final(15 downto 9), "0001101") then                  
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6));    
                    cortex_m0_opcode <= "SUBS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";   
                -------------------------------------------------------------------------------------- -- SUBS <Rdn>,#<imm8> 
                elsif std_match(current_instruction_final(15 downto 11), "00111") then                     
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8));
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "SUBS " & Rd_decode & "," & imm8_decode & "      ";    
                -------------------------------------------------------------------------------------- -- SBCS <Rdn>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "0100000110") then                 
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "SBCS " & Rd_decode & "," & Rm_decode & "       ";   
                -------------------------------------------------------------------------------------- -- RSBS <Rd>,<Rn>,#0 
                elsif std_match(current_instruction_final(15 downto 6), "0100001001") then                 
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "RSBS " & Rd_decode & "," & Rn_decode & "       ";   
                -------------------------------------------------------------------------------------- -- SUB SP,SP,#<imm7> 
                elsif std_match(current_instruction_final(15 downto 7), "101100001") then                 
                    imm8_decode(2) :=   hexcharacter ('0' & current_instruction_final (6 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "SUB SP,SP," & imm8_decode & "    "; 
                    
                -------------------------------------------------------------------------------------- -- MULS <Rdm>,<Rn>,<Rdm>
                elsif std_match(current_instruction_final(15 downto 6), "0100001101") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "MULS " & Rd_decode & "," & Rn_decode & "," & Rd_decode & "    ";  
                -------------------------------------------------------------------------------------- -- CMP <Rn>,<Rm> T1
                elsif std_match(current_instruction_final(15 downto 6), "0100001010") then                
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "CMP  " & Rn_decode & "," & Rm_decode & "       ";   
                -------------------------------------------------------------------------------------- -- CMP <Rn>,<Rm> T2
                elsif std_match(current_instruction_final(15 downto 8), "01000101") then                
                    Rn_decode(2) := hexcharacter (current_instruction_final(7) & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter (current_instruction_final (6 downto 3));
                    cortex_m0_opcode <= "CMP  " & Rn_decode & "," & Rm_decode & "       ";   
                -------------------------------------------------------------------------------------- -- CMN <Rn>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "0100001011") then                
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));
                    cortex_m0_opcode <= "CMN  " & Rn_decode & "," & Rm_decode & "       ";   
                -------------------------------------------------------------------------------------- -- CMP <Rn>,#<imm8> 
                elsif std_match(current_instruction_final(15 downto 11), "00101") then                
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8));
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "CMP  " & Rd_decode & "," & imm8_decode & "      "; 
                -------------------------------------------------------------------------------------- -- ANDS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100000000") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "ANDS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";
                -------------------------------------------------------------------------------------- -- EORS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100000001") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "EORS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";
                -------------------------------------------------------------------------------------- -- ORRS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100001100") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "ORRS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";
                -------------------------------------------------------------------------------------- -- BICS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100001110") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "BICS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";
                -------------------------------------------------------------------------------------- -- MVNS <Rd>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100001111") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "MVNS " & Rd_decode & "," & Rm_decode &  "       "; 
                -------------------------------------------------------------------------------------- -- TST <Rn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100001000") then                
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "TST  " & Rn_decode & "," & Rm_decode &  "       "; 
                -------------------------------------------------------------------------------------- -- LSLS <Rd>,<Rm>,#<imm5>
                elsif std_match(current_instruction_final(15 downto 11), "00000") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));  
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "LSLS " & Rd_decode & "," & Rm_decode & "," & imm8_decode & "   ";  
                -------------------------------------------------------------------------------------- -- LSLS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100000010") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "LSLS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";  
                -------------------------------------------------------------------------------------- -- LSRS <Rd>,<Rm>,#<imm5>
                elsif std_match(current_instruction_final(15 downto 11), "00001") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));  
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "LSRS " & Rd_decode & "," & Rm_decode & "," & imm8_decode & "   ";  
                -------------------------------------------------------------------------------------- -- LSRS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100000011") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "LSRS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";             
                -------------------------------------------------------------------------------------- -- ASRS <Rd>,<Rm>,#<imm5>
                elsif std_match(current_instruction_final(15 downto 11), "00010") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));  
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "ASRS " & Rd_decode & "," & Rm_decode & "," & imm8_decode & "   ";  
                -------------------------------------------------------------------------------------- -- ASRS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100000100") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "ASRS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";             
                -------------------------------------------------------------------------------------- -- RORS <Rdn>,<Rm>
                elsif std_match(current_instruction_final(15 downto 6), "0100000111") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0));
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3));    
                    cortex_m0_opcode <= "RORS " & Rd_decode & "," & Rn_decode & "," & Rm_decode & "    ";
                -------------------------------------------------------------------------------------- -- LDR <Rt>, [<Rn>{,#<imm5>}]
                elsif std_match(current_instruction_final(15 downto 11), "01101") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "LDR  " & Rd_decode & ",[" & Rn_decode & "," & imm8_decode & "] ";  
                -------------------------------------------------------------------------------------- -- LDR <Rt>,[SP{,#<imm8>}]
                elsif std_match(current_instruction_final(15 downto 11), "10011") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8)); -- Rt
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "LDR " & Rd_decode & ",[SP" & "," & imm8_decode & "]  ";  
                -------------------------------------------------------------------------------------- -- LDRH <Rt>, [<Rn>{,#<imm5>}]
                elsif std_match(current_instruction_final(15 downto 11), "10001") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "LDRH " & Rd_decode & ",[" & Rn_decode & "," & imm8_decode & "] ";  
                -------------------------------------------------------------------------------------- -- LDRB <Rt>, [<Rn>{,#<imm5>}]
                elsif std_match(current_instruction_final(15 downto 11), "01111") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "LDRB " & Rd_decode & ",[" & Rn_decode & "," & imm8_decode & "] ";  
                -------------------------------------------------------------------------------------- -- LDR <Rt>,[<Rn>,<Rm>]
                elsif std_match(current_instruction_final(15 downto 9), "0101100") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "LDR  " & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  "; 
                -------------------------------------------------------------------------------------- -- LDRH <Rt>,[<Rn>,<Rm>]
                elsif std_match(current_instruction_final(15 downto 9), "0101101") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "LDRH " & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  ";                  
               ------------------------------------------------------------------------------------- -- LDRSH <Rt>,[<Rn>,<Rm>]
               elsif std_match(current_instruction_final(15 downto 9), "0101111") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "LDRSH" & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  ";                  
                -------------------------------------------------------------------------------------- -- LDRB <Rt>,[<Rn>,<Rm>]
                elsif std_match(current_instruction_final(15 downto 9), "0101110") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "LDRB " & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  ";      
                -------------------------------------------------------------------------------------- -- LDR <Rt>,<label>
                elsif std_match(current_instruction_final(15 downto 11), "01001") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8)); --Rt 
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "LDR  " & Rd_decode & ",[pc," & imm8_decode & "] ";    
                ------------------------------------------------------------------------------------- -- LDM <Rn>!,<registers>
                elsif std_match(current_instruction_final(15 downto 11), "11001") then                
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8)); -- Rn 
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "LDM " & Rd_decode & "!,{" & imm8_decode & "}"  & "    ";   
                 
                -------------------------------------------------------------------------------------- -- STR <Rt>, [<Rn>{,#<imm5>}]
                elsif std_match(current_instruction_final(15 downto 11), "01100") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "STR  " & Rd_decode & ",[" & Rn_decode & "," & imm8_decode & "] ";  
                -------------------------------------------------------------------------------------- -- STRH <Rt>, [<Rn>{,#<imm5>}]
                elsif std_match(current_instruction_final(15 downto 11), "10000") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "STRH " & Rd_decode & ",[" & Rn_decode & "," & imm8_decode & "] ";  
                -------------------------------------------------------------------------------------- -- STRB <Rt>, [<Rn>{,#<imm5>}]
                elsif std_match(current_instruction_final(15 downto 11), "01110") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    imm8_decode(2) :=  hexcharacter ("000" & current_instruction_final (10));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (9 downto 6));  
                    cortex_m0_opcode <= "STRB " & Rd_decode & ",[" & Rn_decode & "," & imm8_decode & "] ";  
                -------------------------------------------------------------------------------------- -- STR <Rt>,[<Rn>,<Rm>]
                elsif std_match(current_instruction_final(15 downto 9), "0101000") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "STR  " & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  ";     
                -------------------------------------------------------------------------------------- -- STRH <Rt>,[<Rn>,<Rm>]
                elsif std_match(current_instruction_final(15 downto 9), "0101001") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "STRH " & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  ";                  
                -------------------------------------------------------------------------------------- -- STRB <Rt>,[<Rn>,<Rm>]
                elsif std_match(current_instruction_final(15 downto 9), "0101010") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rt
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rn 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (8 downto 6)); -- Rm 
                    cortex_m0_opcode <= "STRB " & Rd_decode & ",[" & Rn_decode & "," & Rm_decode & "]  ";     
                -------------------------------------------------------------------------------------- -- STR <Rt>,[SP,#<imm8>]   
                elsif std_match(current_instruction_final(15 downto 11), "10010") then                
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8)); --Rt 
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "STR  " & Rd_decode & ",[sp," & imm8_decode & "] ";      
                ------------------------------------------------------------------------------------- -- STM <Rn>!,<registers>
                elsif std_match(current_instruction_final(15 downto 11), "11000") then                
                    Rn_decode(2) := hexcharacter ('0' & current_instruction_final (10 downto 8)); -- Rn 
                    imm8_decode(2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "STM " & Rn_decode & "!,{" & imm8_decode & "}"  & "    "; 
                ------------------------------------------------------------------------------------- -- PUSH <registers>
                elsif std_match(current_instruction_final(15 downto 9), "1011010") then    
                    LR_PC_decode (2) := hexcharacter ("000" & current_instruction_final (8));            
                    imm8_decode (2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode (3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "PUSH " & "LR=" & LR_PC_decode & ",{" & imm8_decode & "}"  & " ";  
                ------------------------------------------------------------------------------------- -- POP <registers>
                elsif std_match(current_instruction_final(15 downto 9), "1011110") then    
                    LR_PC_decode (2) := hexcharacter ("000" & current_instruction_final (8));            
                    imm8_decode (2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode (3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "POP " & "PC=" & LR_PC_decode & ",{" & imm8_decode & "}"  & "  ";    
                ------------------------------------------------------------------------------------- -- SVC #<imm8>
                elsif std_match(current_instruction_final(15 downto 8), "11011111") then    
                    imm8_decode (2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode (3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "SVC " & ", " & imm8_decode & "        ";                                                                
                ------------------------------------------------------------------------------------- -- B <label>   T1
                elsif std_match(current_instruction_final(15 downto 12), "1101") then    
                    case (current_instruction_final(11 downto 8)) is
                        when EQ => cond_decode := "EQ";
                        when NE => cond_decode := "NE";
                        when CS => cond_decode := "CS"; 
                        when CC => cond_decode := "CC";
                        when MI => cond_decode := "MI";
                        when PL => cond_decode := "PL";
                        when VS => cond_decode := "VS";
                        when VC => cond_decode := "VC";
                        when HI => cond_decode := "HI";
                        when LS => cond_decode := "LS";
                        when GE => cond_decode := "GE";
                        when LT => cond_decode := "LT";
                        when GT => cond_decode := "GT";
                        when LE => cond_decode := "LE";
                        when AL => cond_decode := "AL";
                        when others => cond_decode := "--";
                    end case;         
                    imm8_decode (2) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode (3) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "B" & cond_decode & " ,{" & imm8_decode & "}"  & "       ";
                ------------------------------------------------------------------------------------- -- B <label>   T2
                elsif std_match(current_instruction_final(15 downto 11), "11100") then    
                    imm11_decode (2) :=  hexcharacter ('0' & current_instruction_final (10 downto 8));
                    imm11_decode (3) :=  hexcharacter (current_instruction_final (7 downto 4));
                    imm11_decode (4) :=  hexcharacter (current_instruction_final (3 downto 0));  
                    cortex_m0_opcode <= "B" & " ,{" & imm11_decode & "}"  & "        ";                    
                ------------------------------------------------------------------------------------- -- BL <label>  
    --           elsif std_match(current_instruction_final(15 downto 11), "11110") then    
    --                imm11_decode (2) :=  hexcharacter ('0' & current_instruction_final (10 downto 8));
    --                imm11_decode (3) :=  hexcharacter (current_instruction_final (7 downto 4));
    --                imm11_decode (4) :=  hexcharacter (current_instruction_final (3 downto 0));  
    --                cortex_m0_opcode <= "BL" & " ,{" & imm11_decode & "}"  & "       ";   
                ------------------------------------------------------------------------------------- -- BX Rm  
                elsif std_match(current_instruction_final(15 downto 7), "010001110") then    
                    Rm_decode(2) := hexcharacter (current_instruction_final (6 downto 3)); -- Rm 
                    cortex_m0_opcode <= "BX" & " ," & Rm_decode & "           ";   
                ------------------------------------------------------------------------------------- -- BLX Rm  
                elsif std_match(current_instruction_final(15 downto 7), "010001111") then    
                    Rm_decode(2) := hexcharacter (current_instruction_final (6 downto 3)); -- Rm 
                    cortex_m0_opcode <= "BLX" & " ," & Rm_decode & "          ";                                        
                ------------------------------------------------------------------------------------- -- SXTH <Rd>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "1011001000") then    
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rd 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rm 
                    cortex_m0_opcode <= "SXTH" & " " & Rd_decode & ", " & Rm_decode & "      ";     
                ------------------------------------------------------------------------------------- -- SXTB <Rd>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "1011001001") then    
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rd 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rm 
                    cortex_m0_opcode <= "SXTB" & " " & Rd_decode & ", " & Rm_decode & "      ";  
                ------------------------------------------------------------------------------------- -- REV <Rd>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "1011101000") then    
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rd 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rm 
                    cortex_m0_opcode <= "REV " & " " & Rd_decode & ", " & Rm_decode & "      ";             
                ------------------------------------------------------------------------------------- -- REV16 <Rd>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "1011101001") then    
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rd 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rm 
                    cortex_m0_opcode <= "REV16 " & " " & Rd_decode & ", " & Rm_decode & "    ";             
                ------------------------------------------------------------------------------------- -- REVSH <Rd>,<Rm> 
                elsif std_match(current_instruction_final(15 downto 6), "1011101011") then    
                    Rd_decode(2) := hexcharacter ('0' & current_instruction_final (2 downto 0)); -- Rd 
                    Rm_decode(2) := hexcharacter ('0' & current_instruction_final (5 downto 3)); -- Rm 
                    cortex_m0_opcode <= "REVSH " & " " & Rd_decode & ", " & Rm_decode & "    ";  
                ------------------------------------------------------------------------------------- --  CPS<effect> i 
                elsif std_match(current_instruction_final(15 downto 5), "10110110011") and
                      std_match(current_instruction_final(3 downto 0), "0010") then    
                    imm8_decode(2) :=   hexcharacter (B"0000");
                    imm8_decode(3) :=   hexcharacter (B"000" & current_instruction_final (4));
                    cortex_m0_opcode <= "CPS " & imm8_decode & "          ";         
                ------------------------------------------------------------------------------------- --  BKPT #<imm8>
                elsif std_match(current_instruction_final(15 downto 8), "10111110") then    
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "BKPT " & imm8_decode & "         ";
                ------------------------------------------------------------------------------------- --  SEV
                elsif std_match(current_instruction_final(15 downto 0), "1011111101000000") then    
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "SEV " & imm8_decode & "          ";
                ------------------------------------------------------------------------------------- --  WFI
                elsif std_match(current_instruction_final(15 downto 0), "1011111100110000") then    
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "WFI " & imm8_decode & "          "; 
                ------------------------------------------------------------------------------------- --  YIELD
                elsif std_match(current_instruction_final(15 downto 0), "1011111100010000") then    
                    imm8_decode(2) :=   hexcharacter (current_instruction_final (7 downto 4));
                    imm8_decode(3) :=   hexcharacter (current_instruction_final (3 downto 0));
                    cortex_m0_opcode <= "YIELD " & imm8_decode & "        ";          
              
                end if;
            else -- inst32_detected = true
                -- 32-bit instruction opcode is detected. (HI part)
                cortex_m0_opcode <= "EVAL_32_INSTR    ";  
            end if; -- if (inst32_detected = false)
        end if; -- if (inst32_detected_in_prev_instr = true)
    end if; -- if internal_reset = '1'
    end process;
 
 --synthesis translate on
      
end Behavioral;
